----------------------------------------------------------------------------------
-- Company: McGill University
-- Engineer: Xiangyun Wang
-- 
-- Create Date: 06/18/2021 12:55:30 PM
-- Design Name: BRAM Test
-- Module Name: BRAM_test - Behavioral
-- Project Name: 
-- Target Devices: Arty A7
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
library UNISIM;
use UNISIM.VComponents.all;

entity BRAM_test is
    Port ( 
        DO : out std_logic_vector(7 downto 0);
        ADDR : in std_logic_vector(11 downto 0);
        CLK : in std_ulogic;
        DI : in std_logic_vector(7 downto 0);
        EN : in std_ulogic;
        REGCE : in std_ulogic;
        RST : in std_ulogic;
        WE : in std_logic_vector(0 downto 0));
end BRAM_test;

architecture Behavioral of BRAM_test is

    component BRAM_SINGLE_MACRO is 
        generic (
        --BRAM_SIZE : string := "18Kb";
        --DEVICE : string := "VIRTEX5";
        --DO_REG : integer := 0;
        --INIT : bit_vector := X"000000000000000000";
        --INIT_FILE : string := "NONE";
        --READ_WIDTH : integer := 1;
        --SIM_MODE : string := "SAFE"; -- This parameter is valid only for Virtex5
        --SRVAL : bit_vector := X"000000000000000000";
        --WRITE_MODE : string := "WRITE_FIRST";
        --WRITE_WIDTH : integer := 1;
        
        BRAM_SIZE : string := "36Kb";
        DEVICE : string := "7SERIES";
        DO_REG : integer := 0;
        INIT : bit_vector := X"0000000000";
        INIT_FILE : string := "NONE";
        READ_WIDTH : integer := 8;
        SIM_MODE : string := "SAFE"; -- This parameter is valid only for Virtex5
        SRVAL : bit_vector := X"0000000000";
        WRITE_MODE : string := "WRITE_FIRST";
        WRITE_WIDTH : integer := 8;
        
        --BRAM_SIZE => "36Kb",
        --DEVICE => "7SERIES",
        --DO_REG => 0,
        --INIT => X"0000000000000000",
        --INIT_FILE => "NONE",
        --READ_WIDTH => 16,
        --SIM_MODE => "SAFE", -- This parameter is valid only for Virtex5
        --SRVAL => X"0000000000000000",
        --WRITE_MODE => "WRITE_FIRST",
        --WRITE_WIDTH => 16,
        
        INITP_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INITP_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INITP_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INITP_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INITP_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INITP_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INITP_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INITP_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INITP_08 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INITP_09 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INITP_0A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INITP_0B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INITP_0C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INITP_0D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INITP_0E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INITP_0F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_00 : bit_vector := X"1111111111111111111111111111111111111111111111111111111111111111";
        INIT_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_08 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_09 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_0A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_0B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_0C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_0D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_0E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_0F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_40 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_41 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_42 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_43 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_44 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_45 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_46 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_47 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_48 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_49 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_4A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_4B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_4C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_4D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_4E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_4F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_50 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_51 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_52 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_53 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_54 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_55 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_56 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_57 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_58 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_59 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_5A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_5B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_5C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_5D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_5E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_5F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_60 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_61 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_62 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_63 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_64 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_65 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_66 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_67 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_68 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_69 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_6A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_6B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_6C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_6D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_6E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_6F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_70 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_71 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_72 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_73 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_74 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_75 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_76 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_77 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_78 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_79 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_7A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_7B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_7C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_7D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_7E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
        INIT_7F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
  
      );
    -- ports are unconstrained arrays
    port (
      
        DO : out std_logic_vector(READ_WIDTH-1 downto 0);
        ADDR : in std_logic_vector(11 downto 0);
        CLK : in std_ulogic;
        DI : in std_logic_vector(WRITE_WIDTH-1 downto 0);
        EN : in std_ulogic;
        REGCE : in std_ulogic;
        RST : in std_ulogic;
        WE : in std_logic_vector(0 downto 0)
    
      );
end component;

        --signal DO : std_logic_vector(15 downto 0);
        --signal ADDR : std_logic_vector;
        --signal CLK : std_ulogic;
        --signal DI : std_logic_vector(15 downto 0);
        --signal EN : std_ulogic;
        --signal REGCE : std_ulogic;
        --signal RST : std_ulogic;
        --signal WE : std_logic_vector);

begin

    BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
     generic map(
        BRAM_SIZE => "36Kb",
        DEVICE => "7SERIES",
        DO_REG => 0,
        INIT => X"00000000",
        INIT_FILE => "NONE",
        READ_WIDTH => 8,
        SIM_MODE => "SAFE", -- This parameter is valid only for Virtex5
        SRVAL => X"00000000",
        WRITE_MODE => "WRITE_FIRST",
        WRITE_WIDTH => 8,
        INITP_00  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_01  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_02  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_03  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_04  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_05  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_06  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_07  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_08  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_09  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0A  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0B  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0C  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0D  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0E  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0F  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_00  => X"1111111111111111111111111111111111111111111111111111111111111111",
        INIT_01  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_02  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_03  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_04  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_05  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_06  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_07  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_08  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_09  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0A  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0B  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0C  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0D  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0E  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0F  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_10  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_11  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_12  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_13  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_14  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_15  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_16  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_17  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_18  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_19  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1A  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1B  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1C  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1D  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1E  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1F  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_20  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_21  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_22  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_23  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_24  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_25  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_26  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_27  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_28  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_29  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2A  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2B  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2C  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2D  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2E  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2F  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_30  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_31  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_32  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_33  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_34  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_35  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_36  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_37  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_38  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_39  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3A  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3B  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3C  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3D  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3E  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3F  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_40  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_41  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_42  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_43  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_44  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_45  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_46  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_47  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_48  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_49  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4A  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4B  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4C  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4D  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4E  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4F  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_50  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_51  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_52  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_53  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_54  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_55  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_56  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_57  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_58  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_59  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5A  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5B  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5C  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5D  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5E  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5F  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_60  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_61  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_62  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_63  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_64  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_65  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_66  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_67  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_68  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_69  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6A  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6B  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6C  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6D  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6E  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6F  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_70  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_71  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_72  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_73  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_74  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_75  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_76  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_77  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_78  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_79  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7A  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7B  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7C  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7D  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7E  => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7F  => X"0000000000000000000000000000000000000000000000000000000000000000"
      )
    -- ports are unconstrained arrays
    port map(
      
        DO =>DO,
        ADDR => ADDR,
        CLK => CLK,
        DI => DI,
        EN => EN,
        REGCE => REGCE,
        RST => RST,
        WE => WE
    
      );
      
     -- end of port map
     
     -- customized logic
     -- input signal can be changed
     
end Behavioral;
